
module testbench_4to16;
  reg [3:0]   a;
  reg         en;
  wire [15:0] bcode;

  bindec_4to16 uut(
    .a,
    .en,
    .bcode
  );

  initial begin
    a = 4'b0000;
    en = 'b0;
    # 200;
    a = 4'b0001;
    en = 'b0;
    # 200;
    a = 4'b0010;
    en = 'b0;
    # 200;
    a = 4'b0011;
    en = 'b0;
    # 200;
    a = 4'b0000;
    en = 'b1;
    # 200;
    a = 4'b0001;
    en = 'b1;
    # 200;
    a = 4'b0010;
    en = 'b1;
    # 200;
    a = 4'b0011;
    en = 'b1;
    # 200;
    a = 4'b0100;
    en = 'b0;
    # 200;
    a = 4'b0101;
    en = 'b0;
    # 200;
    a = 4'b0110;
    en = 'b0;
    # 200;
    a = 4'b0111;
    en = 'b0;
    # 200;
    a = 4'b0100;
    en = 'b1;
    # 200;
    a = 4'b0101;
    en = 'b1;
    # 200;
    a = 4'b0110;
    en = 'b1;
    # 200;
    a = 4'b0111;
    en = 'b1;
    # 200;
    a = 4'b1000;
    en = 'b0;
    # 200;
    a = 4'b1001;
    en = 'b0;
    # 200;
    a = 4'b1010;
    en = 'b0;
    # 200;
    a = 4'b1011;
    en = 'b0;
    # 200;
    a = 4'b1000;
    en = 'b1;
    # 200;
    a = 4'b1001;
    en = 'b1;
    # 200;
    a = 4'b1010;
    en = 'b1;
    # 200;
    a = 4'b1011;
    en = 'b1;
    # 200;
    a = 4'b1100;
    en = 'b0;
    # 200;
    a = 4'b1101;
    en = 'b0;
    # 200;
    a = 4'b1110;
    en = 'b0;
    # 200;
    a = 4'b1111;
    en = 'b0;
    # 200;
    a = 4'b1100;
    en = 'b1;
    # 200;
    a = 4'b1101;
    en = 'b1;
    # 200;
    a = 4'b1110;
    en = 'b1;
    # 200;
    a = 4'b1111;
    en = 'b1;
    # 200;
    $stop;
  end
endmodule
